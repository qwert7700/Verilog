

module andGate (
    input wire a,
    input wire b,

    output wire c
);

// changing this file into a verilog file

//This is a file in gitbranch3