

module andGate (
    input wire a,
    input wire b,

    output wire c
);

initial begin 
    a = 0 ;
    b = 0 ;
    c = 0 ;

end 
//Adding changes to a branch

//adding changes to a branch again
//adding another comment 